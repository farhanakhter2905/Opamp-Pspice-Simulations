* F:\Study\2nd year\Analog electronic circuit\New folder\fw.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 20 23:26:08 2021



** Analysis setup **
.tran 0ns 2ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "fw.net"
.INC "fw.als"


.probe


.END
