* F:\Study\2nd year\Analog electronic circuit\lab\l2\sTrigger1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Oct 31 18:58:49 2020



** Analysis setup **
.tran 0ns 30ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "sTrigger1.net"
.INC "sTrigger1.als"


.probe


.END
