* F:\Study\2nd year\Analog electronic circuit\New folder\wien.sch

* Schematics Version 9.1 - Web Update 1
* Sun Mar 21 18:48:45 2021



** Analysis setup **
.tran 1ns 5ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "wien.net"
.INC "wien.als"


.probe


.END
