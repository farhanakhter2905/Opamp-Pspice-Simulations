* F:\Study\2nd year\Analog electronic circuit\lab\LAB 4\6A.sch

* Schematics Version 9.1 - Web Update 1
* Thu Nov 19 00:49:57 2020



** Analysis setup **
.tran 0ns 5ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "6A.net"
.INC "6A.als"


.probe


.END
