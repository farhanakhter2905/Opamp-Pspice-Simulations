* F:\Study\2nd year\Analog electronic circuit\lab\LAB 4\gB.sch

* Schematics Version 9.1 - Web Update 1
* Wed Nov 25 16:14:47 2020



** Analysis setup **
.tran 0ns 2Ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "gB.net"
.INC "gB.als"


.probe


.END
