* F:\Study\2nd year\Analog electronic circuit\lab\LAB 4\pa3.sch

* Schematics Version 9.1 - Web Update 1
* Wed Nov 25 22:16:53 2020



** Analysis setup **
.tran 0ns 2ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "pa3.net"
.INC "pa3.als"


.probe


.END
