* F:\Study\2nd year\Analog electronic circuit\lab\wein2.sch

* Schematics Version 9.1 - Web Update 1
* Sun Mar 21 19:13:57 2021



** Analysis setup **
.tran 1ns 5ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "wein2.net"
.INC "wein2.als"


.probe


.END
