* F:\Study\2nd year\Analog electronic circuit\lab\LAB 4\pa.sch

* Schematics Version 9.1 - Web Update 1
* Wed Nov 25 15:58:43 2020



** Analysis setup **
.tran 0ns 2ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "pa.net"
.INC "pa.als"


.probe


.END
