* F:\Study\2nd year\Analog electronic circuit\lab\l2\oo\Schematic26.sch

* Schematics Version 9.1 - Web Update 1
* Mon Nov 02 14:00:39 2020



** Analysis setup **
.tran 0ns 5ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic26.net"
.INC "Schematic26.als"


.probe


.END
