* F:\Study\2nd year\Analog electronic circuit\lab\l2\SawWave1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Oct 31 20:46:47 2020



** Analysis setup **
.tran 0ns 5ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "SawWave1.net"
.INC "SawWave1.als"


.probe


.END
